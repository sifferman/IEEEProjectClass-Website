
module image (
    input               clk, rst,
    input         [9:0] position_x, position_x_NEXT,
    input         [8:0] position_y, position_y_NEXT,
    input        [31:0] frame,
    output logic  [3:0] r, g, b
);

    // TODO

endmodule
